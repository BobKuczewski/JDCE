5 8 5 0 1
parts.S7400.C74ls279 12 9
parts.input.CPower 7 9
parts.output.CLED_G 13 16
parts.input.CBM_SPDT_I 13 4
parts.input.CBM_SPDT_I 18 4
1 2 2 1 1
3 2 0 6 2
4 2 0 5 2
2 2 0 7 3
1 2 3 3 1
3 3 4 3 1
1 1 3 1 9
3 1 4 1 9
13 15 Q
