3 17 10 0 0
parts.input.CKeyboard 13 12
parts.input.CPower 6 13
parts.output.CBARGRPH8 14 5
1 2 2 1 1
2 1 2 2 1
2 2 2 3 1
2 3 2 4 1
2 4 2 5 1
2 5 2 6 1
2 6 2 7 1
2 7 2 8 1
1 1 0 1 9
0 13 2 9 2
0 14 2 10 2
0 15 2 11 2
0 16 2 12 2
0 17 2 13 2
0 18 2 14 2
0 19 2 15 2
0 20 2 16 2
