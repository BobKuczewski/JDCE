6 12 7 0 0
parts.S7400.C74ls74 9 9
parts.input.CPower 5 9
parts.input.CBT_SPDT_I 9 4
parts.input.CBM_SPDT_I 15 4
parts.input.CBM_SPDT_I 21 9
parts.output.CLED_G 12 16
1 2 2 1 1
2 1 3 1 1
3 1 4 3 1
1 2 5 1 1
1 1 2 3 9
2 3 3 3 9
3 3 4 1 9
2 2 0 2 2
3 2 0 3 2
0 5 5 2 3
4 2 0 1 5
0 6 0 4 11
