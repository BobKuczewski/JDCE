; Header Line:  NumParts, NumWires, NumNets, NumProbes, NumLabels

6 44 24 24 2

; Parts List:   Package.Class, LocationX, LocationY, optional parameters

parts.cdp1800.CCDP1802BC 20 18  ; 1802 located at grid point (20,18)
parts.rom.C2708 28 32 Blink_Q   ; This is a ROM from file "Blink_Q.rom"
parts.input.CClock 25 12        ; Clock chip
parts.input.CPower 14 28        ; Power for the circuit
parts.S7400.C74ls91 15 12       ; Shift register to provide delayed reset
parts.output.CLED_R 23 29       ; Q Output LED

; Wires List:   PartNum,PinNum, PartNum,PinNum, Color

1 17 0 8 2
0 9 1 16 2
1 15 0 10 2
1 13 0 12 2
1 11 0 13 2
1 10 0 14 2
1 9 0 15 2
1 20 0 7 11
0 25 1 8 5
0 26 1 7 5
0 27 1 6 5
1 5 0 28 5
0 29 1 4 5
1 3 0 30 5
0 31 1 2 5
2 1 0 1 5    ; 1802's Pin1 (CLK) from Clock's Pin1
3 2 1 19 1
1 19 1 22 1
1 22 1 23 1
1 19 1 18 1
1 18 1 12 1
3 2 0 20 1
3 1 0 2 9
0 35 0 36 9
3 1 0 40 9
0 32 1 1 5
0 11 1 14 2
4 9 2 2 3
3 1 4 12 9
3 2 4 10 1
4 12 4 11 9
0 3 4 13 3
4 5 4 11 9
3 1 1 24 9
0 4 5 2 11   ; 1802's Pin4 (Q) to LED's Pin2
5 1 3 2 1
0 36 0 37 9
0 37 0 38 9
0 38 3 1 9
0 16 4 11 9
0 16 0 24 9
0 24 0 23 9
0 23 0 22 9
0 22 0 21 9

; Probes List:  PartNum, PinNum, DisplayName

0 3 /CLR
0 1 CLK
0 34 TPA
0 33 TPB
0 6 SC0
0 7 /MRD
0 35 /MWR
0 32 A7
0 31 A6
0 30 A5
0 29 A4
0 28 A3
0 27 A2
0 26 A1
0 25 A0
0 8 D7
0 9 D6
0 10 D5
0 11 D4
0 12 D3
0 13 D2
0 14 D1
0 15 D0
0 4 Q

; Labels List:  LocationX, LocationY, Text

12 36 Simple 1802
12 38 with 256 byte ROM
