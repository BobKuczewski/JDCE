22 56 22 0 0
parts.S7400.C74ls181 19 24
parts.input.CPower 12 25
parts.input.CBT_SPDT_I 19 18
parts.input.CBT_SPDT_I 22 18
parts.input.CBT_SPDT_I 25 18
parts.input.CBT_SPDT_I 28 18
parts.input.CBT_SPDT_I 19 12
parts.input.CBT_SPDT_I 22 12
parts.input.CBT_SPDT_I 25 12
parts.input.CBT_SPDT_I 28 12
parts.output.CLED_G 19 35
parts.output.CLED_G 22 35
parts.output.CLED_G 25 35
parts.output.CLED_G 28 35
parts.input.CBT_SPDT_I 34 18
parts.input.CBT_SPDT_I 37 18
parts.input.CBT_SPDT_I 40 18
parts.input.CBT_SPDT_I 43 18
parts.input.CBT_SPDT_I 35 25
parts.input.CBT_SPDT_I 34 12
parts.input.CBT_SPDT_I 40 12
parts.input.CBT_SPDT_I 43 12
1 2 2 1 1
2 1 3 1 1
3 1 4 1 1
4 1 5 1 1
1 2 6 1 1
6 1 7 1 1
7 1 8 1 1
8 1 9 1 1
1 1 2 3 9
2 3 3 3 9
3 3 4 3 9
4 3 5 3 9
1 1 6 3 9
6 3 7 3 9
7 3 8 3 9
8 3 9 3 9
1 2 10 1 1
10 1 11 1 1
11 1 12 1 1
12 1 13 1 1
5 1 14 1 1
14 1 15 1 1
15 1 16 1 1
16 1 17 1 1
5 3 14 3 9
14 3 15 3 9
15 3 16 3 9
16 3 17 3 9
5 2 0 2 2
9 2 0 1 2
4 2 0 23 2
8 2 0 22 2
3 2 0 21 2
7 2 0 20 2
2 2 0 19 2
6 2 0 18 2
14 2 0 3 6
15 2 0 4 6
16 2 0 5 6
17 2 0 6 6
0 9 13 2 3
0 10 12 2 3
0 11 11 2 3
0 13 10 2 3
5 1 18 1 1
5 3 18 3 9
18 2 0 8 5
9 1 19 1 1
9 3 19 3 9
19 2 0 7 2
19 1 20 1 1
20 1 21 1 1
19 3 20 3 9
20 3 21 3 9
20 2 0 15 5
21 2 0 17 5
