15 47 21 0 0
parts.rom.C2708 23 22 test
parts.output.CTIL311 23 15
parts.output.CTIL311 31 15
parts.input.CPower 12 23
parts.input.CBT_SPDT_I 12 35
parts.input.CBT_SPDT_I 15 35
parts.input.CBT_SPDT_I 20 35
parts.input.CBT_SPDT_I 23 35
parts.input.CBT_SPDT_I 26 35
parts.input.CBT_SPDT_I 29 35
parts.input.CBT_SPDT_I 33 35
parts.input.CBT_SPDT_I 36 35
parts.input.CBT_SPDT_I 39 35
parts.input.CBT_SPDT_I 42 35
parts.input.CBT_SPDT_I 40 23
3 2 1 5 1
1 5 1 8 1
1 8 2 5 1
2 5 2 8 1
2 3 0 9 5
2 2 0 10 5
2 13 0 11 5
2 12 0 13 5
1 3 0 14 5
1 2 0 15 5
1 13 0 16 5
1 12 0 17 5
3 1 1 1 9
1 1 2 1 9
3 2 4 1 1
4 1 5 1 1
5 1 6 1 1
6 1 7 1 1
7 1 8 1 1
8 1 9 1 1
9 1 10 1 1
10 1 11 1 1
11 1 12 1 1
12 1 13 1 1
3 1 4 3 9
4 3 5 3 9
5 3 6 3 9
6 3 7 3 9
7 3 8 3 9
8 3 9 3 9
9 3 10 3 9
10 3 11 3 9
11 3 12 3 9
12 3 13 3 9
13 1 14 1 1
14 3 13 3 9
14 2 0 20 11
13 2 0 8 2
12 2 0 7 2
11 2 0 6 2
10 2 0 5 2
9 2 0 4 2
8 2 0 3 2
7 2 0 2 2
6 2 0 1 2
5 2 0 23 2
4 2 0 22 2
