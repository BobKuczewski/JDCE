32 188 63 0 0
parts.cpu.C8080A 25 28
parts.output.CTIL311 25 44
parts.output.CTIL311 30 44
parts.output.CTIL311 35 44
parts.output.CTIL311 40 44
parts.input.CPower 6 29
parts.output.CTIL311 50 44
parts.output.CTIL311 55 44
parts.input.CClock 13 29
parts.S7400.C74265 13 36
parts.rom.C2764 25 17 boot8080
parts.ram.CCDM6264 25 6
parts.S7400.C74ls138 13 19
parts.input.CBT_SPDT_I 7 7
parts.input.CBM_SPDT_I 12 7
parts.input.CBT_SPDT_I 17 7
parts.S7400.C74ls04 50 22
parts.S7400.C74ls32 62 22
parts.S7400.C74ls138 50 29
parts.S7400.C74ls373 62 29
parts.S7400.C74ls244 54 14
parts.input.CBT_SPDT_I 49 6
parts.input.CBT_SPDT_I 52 6
parts.input.CBT_SPDT_I 55 6
parts.input.CBT_SPDT_I 46 6
parts.input.CBT_SPDT_I 59 6
parts.input.CBT_SPDT_I 62 6
parts.input.CBT_SPDT_I 65 6
parts.input.CBT_SPDT_I 68 6
parts.output.CBARGRPH8 63 40
parts.output.CLED_R 44 21
parts.output.CLED_R 44 15
5 2 1 5 1
1 5 1 8 1
1 8 2 5 1
2 5 2 8 1
2 8 3 5 1
3 5 3 8 1
3 8 4 5 1
4 5 4 8 1
5 1 1 1 9
1 1 2 1 9
2 1 3 1 9
3 1 4 1 9
0 25 4 3 11
0 26 4 2 11
0 27 4 13 11
0 29 4 12 11
0 30 3 3 11
0 32 3 13 11
0 33 3 12 11
0 34 2 3 11
0 35 2 2 11
0 1 2 13 11
0 40 2 12 11
0 37 1 3 11
0 38 1 2 11
0 39 1 13 11
0 36 1 12 11
4 8 6 8 1
6 8 7 8 1
0 10 7 3 2
0 9 7 2 2
0 8 7 13 2
0 7 7 12 2
0 3 6 3 2
0 4 6 2 2
0 5 6 13 2
0 6 6 12 2
8 2 9 1 5
9 2 0 22 5
9 3 0 15 5
4 1 6 1 9
6 1 7 1 9
5 2 10 20 1
5 2 12 4 1
12 4 12 5 1
12 5 11 22 1
5 1 12 6 9
12 6 11 26 9
13 2 0 13 5
14 2 0 12 5
15 2 0 23 5
0 3 10 16 2
10 16 11 16 2
0 4 10 17 2
10 17 11 17 2
0 5 10 18 2
10 18 11 18 2
0 6 10 19 2
10 19 11 19 2
0 7 10 15 2
10 15 11 15 2
0 8 10 13 2
10 13 11 13 2
0 9 10 12 2
10 12 11 12 2
0 10 10 11 2
10 11 11 11 2
0 25 10 10 11
10 10 11 10 11
0 26 10 9 11
10 9 11 9 11
4 13 0 27 11
0 27 10 8 11
10 8 11 8 11
4 12 0 28 11
0 28 10 7 11
10 7 11 7 11
0 30 10 6 11
10 6 11 6 11
3 2 0 31 11
0 31 10 5 11
10 5 11 5 11
0 32 10 4 11
10 4 11 4 11
0 33 10 3 11
10 3 11 3 11
0 34 10 25 11
10 25 11 25 11
0 35 10 24 11
10 24 11 24 11
0 1 10 21 11
10 21 11 21 11
0 40 10 23 11
10 23 11 23 11
0 37 10 2 11
10 2 11 2 11
0 38 12 1 11
0 39 12 2 11
0 36 12 3 11
12 15 10 22 5
12 14 11 20 5
11 27 0 18 5
5 1 13 3 9
13 3 14 3 9
14 3 15 1 9
5 2 13 1 1
13 1 14 1 1
14 1 15 3 1
16 1 17 6 4
16 2 19 11 5
0 17 16 9 5
16 8 17 13 4
0 25 18 1 11
0 26 18 2 11
0 27 18 3 11
12 7 18 4 5
18 4 18 5 5
5 1 18 6 9
18 13 17 12 5
18 14 17 5 4
18 15 17 1 5
17 3 6 5 4
6 5 7 5 4
0 18 17 2 5
17 2 17 4 5
17 11 20 19 5
20 19 20 1 5
15 3 24 1 1
24 1 21 1 1
21 1 22 1 1
22 1 23 1 1
23 1 25 1 1
25 1 26 1 1
26 1 27 1 1
27 1 28 1 1
15 1 24 3 9
24 3 21 3 9
21 3 22 3 9
22 3 23 3 9
23 3 25 3 9
25 3 26 3 9
26 3 27 3 9
27 3 28 3 9
28 2 20 2 6
27 2 20 4 6
26 2 20 6 6
25 2 20 8 6
23 2 20 11 6
22 2 20 13 6
21 2 20 15 6
24 2 20 17 6
6 3 19 13 2
19 13 20 9 2
6 2 19 14 2
19 14 20 7 2
6 13 19 17 2
19 17 20 5 2
6 12 19 18 2
19 18 20 3 2
7 3 19 3 2
19 3 20 18 2
7 2 19 4 2
19 4 20 16 2
7 13 19 7 2
19 7 20 14 2
7 12 19 8 2
19 8 20 12 2
7 8 29 1 1
29 1 29 2 1
29 2 29 3 1
29 3 29 4 1
29 4 29 5 1
29 5 29 6 1
29 6 29 7 1
29 7 29 8 1
29 9 19 2 6
29 10 19 5 6
29 11 19 6 6
29 12 19 9 6
29 13 19 12 6
29 14 19 15 6
29 15 19 16 6
29 16 19 19 6
7 8 19 1 1
24 1 31 1 1
31 1 30 1 1
31 2 0 21 5
30 2 0 24 5
