9 23 9 0 0
parts.input.CPower 9 11
parts.input.CBT_SPDT_I 17 19
parts.input.CBT_SPDT_I 21 19
parts.input.CBT_SPDT_I 25 19
parts.input.CBT_SPDT_I 29 19
parts.input.CBT_SPDT_I 15 11
parts.output.CTIL311 21 15
parts.input.CBT_SPDT_I 29 14
parts.input.CBT_SPDT_I 33 14
0 2 5 1 1
0 2 1 1 1
1 1 2 1 1
2 1 3 1 1
3 1 4 1 1
5 1 6 5 1
6 5 6 8 1
0 1 5 3 9
0 1 1 3 9
1 3 2 3 9
2 3 3 3 9
3 3 4 3 9
5 2 6 1 2
4 2 6 3 2
3 2 6 2 2
2 2 6 13 2
1 2 6 12 2
7 2 6 4 2
8 2 6 10 2
4 1 8 3 1
8 3 7 3 1
4 3 8 1 9
8 1 7 1 9
