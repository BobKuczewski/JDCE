6 12 6 0 4
parts.S7400.C74ls00 16 16
parts.input.CPower 10 16
parts.output.CLED_R 17 10
parts.output.CLED_G 21 10
parts.input.CBM_SPDT_I 16 23
parts.input.CBM_SPDT_I 22 23
1 2 2 1 1
2 1 3 1 1
4 2 0 1 2
5 2 0 5 2
0 3 2 2 11
0 6 3 2 11
0 3 0 4 11
0 6 0 2 11
1 2 4 3 1
4 3 5 3 1
1 1 4 1 9
4 1 5 1 9
20 8 Q
16 8 /Q
21 21 Set
14 21 Reset
