11 23 11 0 1
parts.S7400.C74ls175 13 12
parts.input.CPower 8 12
parts.input.CBT_SPDT_I 11 6
parts.input.CBT_SPDT_I 15 6
parts.input.CBT_SPDT_I 19 6
parts.input.CBT_SPDT_I 23 6
parts.output.CLED_G 15 19
parts.output.CLED_G 18 19
parts.output.CLED_G 21 19
parts.output.CLED_G 12 19
parts.input.CBM_SPDT_I 27 12
1 2 2 1 1
2 1 3 1 1
3 1 4 1 1
4 1 5 1 1
1 2 9 1 1
9 1 6 1 1
6 1 7 1 1
7 1 8 1 1
5 1 10 1 1
1 1 2 3 9
2 3 3 3 9
3 3 4 3 9
4 3 5 3 9
5 3 10 3 9
5 2 0 4 2
4 2 0 5 2
3 2 0 12 2
2 2 0 13 2
0 2 8 2 3
0 7 7 2 3
0 10 6 2 3
0 15 9 2 3
0 9 10 2 5
26 11 Write
