8 24 14 0 0
parts.cpu.CZ86E08 13 14 etest
parts.output.CTIL311 13 9
parts.output.CTIL311 19 9
parts.input.CPower 6 14
parts.pic.C24LC256 14 22 test
parts.input.CClock 25 14
parts.output.CLED_R 26 7
parts.output.CLED_R 29 7
5 1 0 7 11
0 15 4 5 2
0 15 2 3 2
0 16 2 2 2
0 17 2 13 2
0 18 2 12 2
0 1 1 3 2
0 2 1 2 2
0 3 1 13 2
0 4 1 12 2
0 11 4 6 13
3 2 4 1 1
4 1 4 2 1
4 2 4 3 1
0 12 2 5 13
0 13 1 5 13
3 2 1 8 1
1 8 2 8 1
3 1 1 1 12
1 1 2 1 12
2 8 6 1 1
6 1 7 1 1
0 12 7 2 13
0 13 6 2 13
