5 9 5 0 3
parts.S7400.C74ls74 11 10
parts.input.CPower 6 10
parts.input.CBM_SPDT_I 14 4
parts.input.CBM_SPDT_I 24 10
parts.output.CLED_G 14 17
1 2 2 1 1
2 1 3 3 1
1 1 2 3 9
2 3 3 1 9
1 2 4 1 1
2 3 0 2 9
2 2 0 3 2
0 5 4 2 3
3 2 0 1 5
23 9 Reset
13 3 Pulse
12 16 Output
