19 60 21 0 0
parts.input.CPower 7 15
parts.ram.C2114 14 15
parts.output.CBARGRPH4 15 8
parts.input.CBT_SPDT_I 10 25
parts.input.CBT_SPDT_I 13 25
parts.input.CBT_SPDT_I 16 25
parts.input.CBT_SPDT_I 19 25
parts.input.CBT_SPDT_I 22 25
parts.input.CBT_SPDT_I 26 25
parts.input.CBT_SPDT_I 29 25
parts.input.CBT_SPDT_I 32 25
parts.input.CBT_SPDT_I 35 25
parts.input.CBT_SPDT_I 38 25
parts.S7400.C74ls244 14 34
parts.input.CBT_SPDT_I 12 41
parts.input.CBT_SPDT_I 15 41
parts.input.CBT_SPDT_I 18 41
parts.input.CBT_SPDT_I 21 41
parts.input.CBM_SPDT_I 32 14
0 2 2 1 1
2 1 2 2 1
2 2 2 3 1
2 3 2 4 1
0 2 3 1 1
3 1 4 1 1
4 1 5 1 1
5 1 6 1 1
6 1 7 1 1
7 1 8 1 1
8 1 9 1 1
9 1 10 1 1
10 1 11 1 1
11 1 12 1 1
0 1 3 3 9
3 3 4 3 9
4 3 5 3 9
5 3 6 3 9
6 3 7 3 9
7 3 8 3 9
8 3 9 3 9
9 3 10 3 9
10 3 11 3 9
11 3 12 3 9
12 2 1 5 5
11 2 1 6 5
10 2 1 7 5
9 2 1 4 5
8 2 1 3 5
7 2 1 2 5
6 2 1 1 5
5 2 1 17 5
4 2 1 16 5
3 2 1 15 5
1 11 2 8 2
1 12 2 7 2
1 13 2 6 2
1 14 2 5 2
0 2 14 1 1
14 1 15 1 1
15 1 16 1 1
16 1 17 1 1
0 1 14 3 9
14 3 15 3 9
15 3 16 3 9
16 3 17 3 9
17 2 13 2 6
16 2 13 4 6
15 2 13 6 6
14 2 13 8 6
13 18 2 5 2
13 16 2 6 2
13 14 2 7 2
13 12 2 8 2
2 4 1 8 1
18 3 12 1 1
18 1 12 3 9
18 2 1 10 11
18 2 13 1 11
13 1 13 19 11
