20 90 59 0 5
parts.S7400.C74ls47 9 16
parts.S7400.C74ls47 18 16
parts.S7400.C74ls47 27 16
parts.S7400.C74ls47 36 16
parts.output.CMAN10A 11 12
parts.output.CMAN10A 20 12
parts.output.CMAN10A 29 12
parts.output.CMAN10A 38 12
parts.S7400.C74ls160 9 24
parts.S7400.C74ls160 18 24
parts.S7400.C74ls160 27 24
parts.S7400.C74ls160 36 24
parts.input.CClock 36 32
parts.S7400.C74ls367 36 40
parts.input.CPower 4 34
parts.input.CBM_SPDT_I 12 40
parts.input.CBT_SPDT_I 21 40
parts.input.CBM_SPDT_I 21 32
parts.input.CBT_SPDT_I 30 32
parts.input.CBM_SPDT_I 30 40
4 7 0 9 4
5 7 1 9 4
6 7 2 9 4
7 7 3 9 4
4 2 0 15 4
5 2 1 15 4
6 2 2 15 4
7 2 3 15 4
4 1 0 13 4
5 1 1 13 4
6 1 2 13 4
7 1 3 13 4
4 13 0 12 4
5 13 1 12 4
6 13 2 12 4
7 13 3 12 4
4 11 0 14 4
5 11 1 14 4
6 11 2 14 4
7 11 3 14 4
4 10 0 11 4
5 10 1 11 4
6 10 2 11 4
7 10 3 11 4
4 8 0 10 4
5 8 1 10 4
6 8 2 10 4
7 8 3 10 4
14 1 4 14 9
4 14 5 14 9
5 14 6 14 9
6 14 7 14 9
0 1 8 13 2
1 1 9 13 2
2 1 10 13 2
3 1 11 13 2
0 2 8 12 2
1 2 9 12 2
2 2 10 12 2
3 2 11 12 2
0 3 15 2 3
1 3 15 2 3
2 3 15 2 3
3 3 15 2 3
14 1 15 1 9
14 2 15 3 1
0 4 13 9 5
0 4 1 5 3
1 4 2 5 3
1 4 13 7 5
2 4 13 5 5
3 4 13 3 5
0 5 16 2 3
15 1 16 1 9
15 3 16 3 1
0 6 8 11 2
1 6 9 11 2
2 6 10 11 2
3 6 11 11 2
0 7 8 14 2
1 7 9 14 2
2 7 10 14 2
3 7 11 14 2
14 1 17 1 9
14 2 17 3 1
17 2 8 1 2
17 2 9 1 2
17 2 10 1 2
17 2 11 1 2
8 2 9 15 11
9 2 10 15 11
10 2 11 15 11
11 2 12 1 11
18 2 11 10 5
11 10 11 7 5
18 2 10 10 5
10 10 10 7 5
18 2 9 10 5
9 10 9 7 5
18 2 8 10 5
8 10 8 7 5
17 3 18 1 1
17 1 18 3 9
16 3 13 10 1
13 10 13 6 1
13 6 13 4 1
13 4 13 2 1
19 2 13 1 5
16 1 19 1 9
16 3 19 3 1
11 44 TEST
19 44 LZBLANK
20 36 CLR
29 36 COUNT
29 44 BLANK
