6 37 13 19 0
parts.cdp1800.CCDP1802BC 20 18
parts.input.CClock 25 12
parts.input.CPower 14 28
parts.S7400.C74ls91 15 12
parts.cd4000.CCD4011 36 12
parts.output.CLED_R 28 28
1 1 0 1 5
2 2 0 20 1
2 1 0 2 9
0 35 0 36 9
2 1 0 40 9
3 9 1 2 3
2 1 3 12 9
2 2 3 10 1
3 12 3 11 9
0 3 3 13 3
3 5 3 11 9
0 25 4 12 5
0 26 4 13 2
4 13 4 1 2
4 13 4 2 2
4 11 0 11 11
0 11 0 10 11
4 3 0 14 3
0 14 0 12 3
0 12 0 9 3
0 8 2 2 1
0 13 2 2 1
4 12 4 9 5
4 3 4 8 3
4 10 4 6 6
4 10 4 5 6
4 4 0 15 6
0 4 5 2 5
5 1 2 2 1
3 11 0 16 9
0 16 0 24 9
0 24 0 23 9
0 23 0 22 9
0 22 0 21 9
0 36 0 37 9
0 37 0 38 9
0 38 2 1 9
0 3 /CLR
0 1 CLK
0 34 TPA
0 33 TPB
0 6 SC0
0 7 /MRD
0 35 /MWR
0 27 A2
0 26 A1
0 25 A0
0 8 D7
0 9 D6
0 10 D5
0 11 D4
0 12 D3
0 13 D2
0 14 D1
0 15 D0
0 4 Q
