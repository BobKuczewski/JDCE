15 101 38 0 2
parts.cdp1800.CCDP1802BC 14 20
parts.rom.C2708 38 20 boot1802
parts.ram.CCDM6116A 53 20
parts.output.CTIL311 14 43
parts.output.CTIL311 19 43
parts.output.CTIL311 24 43
parts.output.CTIL311 29 43
parts.output.CTIL311 37 43
parts.output.CTIL311 42 43
parts.input.CPower 4 22
parts.input.CClock 14 13
parts.S7400.C74ls373 19 30
parts.S7400.C74ls04 31 13
parts.input.CBT_SPDT_I 9 22
parts.S7400.C74ls00 42 13
9 2 3 5 1
3 5 3 8 1
3 8 4 5 1
4 5 4 8 1
9 1 3 1 9
3 1 4 1 9
4 1 5 1 9
5 1 6 1 9
6 1 7 1 9
7 1 8 1 9
6 8 7 8 1
7 8 8 8 1
0 25 6 3 11
0 26 6 2 11
0 27 6 13 11
0 28 6 12 11
0 29 5 3 11
0 30 5 2 11
0 31 5 13 11
0 32 5 12 11
10 1 0 1 5
0 15 8 3 2
0 14 8 2 2
0 13 8 13 2
0 12 8 12 2
0 11 7 3 2
0 10 7 2 2
0 9 7 13 2
0 8 7 12 2
8 3 1 9 2
8 2 1 10 2
8 13 1 11 2
8 12 1 13 2
7 3 1 14 2
7 2 1 15 2
7 13 1 16 2
7 12 1 17 2
8 3 2 9 2
8 2 2 10 2
8 13 2 11 2
8 12 2 13 2
7 3 2 14 2
7 2 2 15 2
7 13 2 16 2
7 12 2 17 2
0 25 11 3 11
0 26 11 4 11
0 27 11 7 11
0 28 11 8 11
0 29 11 13 11
0 30 11 14 11
0 31 11 17 11
0 32 11 18 11
11 2 4 3 11
11 5 4 2 11
11 6 4 13 11
11 9 4 12 11
11 12 3 3 11
11 15 3 2 11
11 16 3 13 11
11 19 3 12 11
6 3 1 8 11
6 2 1 7 11
6 13 1 6 11
6 12 1 5 11
5 3 1 4 11
5 2 1 3 11
5 13 1 2 11
5 12 1 1 11
3 12 1 20 11
9 2 13 1 1
9 1 13 3 9
13 2 0 3 5
9 2 11 1 1
0 34 11 11 5
0 22 12 1 5
7 5 8 5 5
4 8 5 8 1
5 8 6 8 1
0 33 12 3 5
12 4 5 5 5
5 5 6 5 5
4 3 1 23 11
4 2 1 22 11
6 3 2 8 11
6 2 2 7 11
6 13 2 6 11
6 12 2 5 11
5 3 2 4 11
5 2 2 3 11
5 13 2 2 11
5 12 2 1 11
4 3 2 23 11
4 2 2 22 11
2 21 0 35 5
2 20 0 7 5
3 12 12 5 11
12 6 2 18 11
7 5 14 3 5
14 2 0 33 5
0 19 14 1 5
8 26 Run
7 21 Reset
