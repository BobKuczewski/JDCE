8 22 10 0 0
parts.pld.C5C031 16 8 ior
parts.output.CBARGRPH4 17 2
parts.input.CPower 7 8
parts.input.CBT_SPDT_I 12 16
parts.input.CBT_SPDT_I 15 16
parts.input.CBT_SPDT_I 18 16
parts.input.CBT_SPDT_I 21 16
parts.input.CBT_SPDT_I 26 16
2 2 1 1 1
1 1 1 2 1
1 2 1 3 1
1 3 1 4 1
2 2 3 1 1
3 1 4 1 1
4 1 5 1 1
5 1 6 1 1
6 1 7 1 1
2 1 3 3 9
3 3 4 3 9
4 3 5 3 9
5 3 6 3 9
6 3 7 3 9
3 2 0 1 2
4 2 0 2 2
5 2 0 3 2
6 2 0 4 2
7 2 0 5 2
0 19 1 5 6
0 18 1 6 6
0 17 1 7 6
