22 60 30 0 0
parts.S7400.C74ls138 12 14
parts.S7400.C74ls138 36 14
parts.output.CLED_R 11 21
parts.output.CLED_R 11 26
parts.output.CLED_R 11 31
parts.output.CLED_R 16 26
parts.output.CLED_R 21 26
parts.output.CLED_R 21 21
parts.output.CLED_R 21 31
parts.S7400.C74ls69 25 21
parts.input.CClock 25 28
parts.S7400.C74ls10 12 36
parts.input.CBT_DPDT_I 26 14
parts.S7400.C74ls10 36 36
parts.output.CLED_R 35 21
parts.output.CLED_R 35 26
parts.output.CLED_R 35 31
parts.output.CLED_R 40 26
parts.output.CLED_R 45 26
parts.output.CLED_R 45 21
parts.output.CLED_R 45 31
parts.input.CPower 4 24
21 2 2 1 1
2 1 7 1 1
21 2 3 1 1
3 1 5 1 1
5 1 6 1 1
6 1 15 1 1
15 1 17 1 1
17 1 18 1 1
17 1 19 1 1
17 1 14 1 1
17 1 20 1 1
17 1 16 1 1
21 2 0 4 1
0 4 0 5 1
0 5 1 4 1
1 4 1 5 1
21 2 4 1 1
4 1 8 1 1
21 1 0 6 9
0 6 1 6 9
2 2 8 2 2
8 2 11 6 2
14 2 20 2 2
20 2 13 6 2
5 2 11 8 2
17 2 13 8 2
4 2 7 2 2
7 2 0 15 2
0 15 11 9 2
16 2 19 2 2
19 2 1 15 2
1 15 13 9 2
3 2 6 2 2
3 2 11 12 2
15 2 18 2 2
15 2 13 12 2
11 3 0 12 2
13 3 1 12 2
11 4 0 11 2
11 4 11 11 2
13 4 1 11 2
13 4 13 11 2
11 5 0 10 2
0 10 11 13 2
13 5 1 10 2
1 10 13 13 2
11 10 0 13 2
13 10 1 13 2
12 2 9 15 11
12 5 9 9 11
9 2 1 1 5
9 3 1 3 5
9 4 1 9 5
9 5 0 3 5
9 7 0 1 5
9 10 0 2 5
9 11 0 9 5
9 13 1 2 5
12 3 10 2 11
10 1 12 6 11
