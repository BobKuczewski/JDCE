8 54 23 0 0
parts.S7400.C74ls138 23 18
parts.S7400.C74ls238 44 18
parts.input.CPower 37 18
parts.input.CBT_SPDT_I 34 25
parts.input.CBT_SPDT_I 37 25
parts.input.CBT_SPDT_I 40 25
parts.output.CBARGRPH8 23 28
parts.output.CBARGRPH8 44 28
2 1 0 16 9
2 1 1 16 9
2 2 0 8 1
2 2 1 8 1
2 1 0 6 9
2 1 1 6 9
2 2 0 5 1
2 2 0 4 1
2 2 1 5 1
2 2 1 4 1
5 2 0 1 2
4 2 0 2 2
3 2 0 3 2
2 2 6 8 1
6 8 6 7 1
6 7 6 6 1
6 6 6 5 1
6 5 6 4 1
6 4 6 3 1
6 3 6 2 1
6 2 6 1 1
0 15 6 9 2
0 14 6 10 2
0 13 6 11 2
0 12 6 12 2
0 11 6 13 2
0 10 6 14 2
0 9 6 15 2
0 7 6 16 2
2 2 7 1 1
7 1 7 2 1
7 2 7 3 1
7 3 7 4 1
7 4 7 5 1
7 5 7 6 1
7 6 7 7 1
7 7 7 8 1
1 15 7 9 2
1 14 7 10 2
1 13 7 11 2
1 12 7 12 2
1 11 7 13 2
1 10 7 14 2
1 9 7 15 2
1 7 7 16 2
5 3 4 3 9
3 3 4 3 9
2 1 5 3 9
4 1 5 1 1
3 1 4 1 1
3 1 2 2 1
3 2 1 3 2
4 2 1 2 2
5 2 1 1 2
